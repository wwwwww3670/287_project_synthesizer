library ieee;
use ieee.std_logic_1164.all;

package sine_package is

  constant max_table_value: integer := 32764;
  subtype table_value_type is integer range -max_table_value to max_table_value;

  constant max_table_index: integer := 127;
  subtype table_index_type is integer range 0 to max_table_index;

  subtype sine_vector_type is std_logic_vector( 15 downto 0 );

  function get_table_value (table_index: table_index_type) return table_value_type;

end;

package body sine_package is

  function get_table_value (table_index: table_index_type) return table_value_type is
    variable table_value: table_value_type;
  begin
    case table_index is
      when 0 =>
        table_value := 0;
      when 1 =>
        table_value := 402;
      when 2 =>
        table_value := 804;
      when 3 =>
        table_value := 1206;
      when 4 =>
        table_value := 1607;
      when 5 =>
        table_value := 2009;
      when 6 =>
        table_value := 2410;
      when 7 =>
        table_value := 2811;
      when 8 =>
        table_value := 3211;
      when 9 =>
        table_value := 3611;
      when 10 =>
        table_value := 4011;
      when 11 =>
        table_value := 4409;
      when 12 =>
        table_value := 4807;
      when 13 =>
        table_value := 5205;
      when 14 =>
        table_value := 5601;
      when 15 =>
        table_value := 5997;
      when 16 =>
        table_value := 6392;
      when 17 =>
        table_value := 6786;
      when 18 =>
        table_value := 7179;
      when 19 =>
        table_value := 7571;
      when 20 =>
        table_value := 7961;
      when 21 =>
        table_value := 2351;
      when 22 =>
        table_value := 8739;
      when 23 =>
        table_value := 9126;
      when 24 =>
        table_value := 9511;
      when 25 =>
        table_value := 9895;
      when 26 =>
        table_value := 10278;
      when 27 =>
        table_value := 10659;
      when 28 =>
        table_value := 11038;
      when 29 =>
        table_value := 11416;
      when 30 =>
        table_value := 11792;
      when 31 =>
        table_value := 12166;
      when 32 =>
        table_value := 12539;
      when 33 =>
        table_value := 12909;
      when 34 =>
        table_value := 13278;
      when 35 =>
        table_value := 13645;
      when 36 =>
        table_value := 14009;
      when 37 =>
        table_value := 14372;
      when 38 =>
        table_value := 14732;
      when 39 =>
        table_value := 15090;
      when 40 =>
        table_value := 15446;
      when 41 =>
        table_value := 15799;
      when 42 =>
        table_value := 16150;
      when 43 =>
        table_value := 16499;
      when 44 =>
        table_value := 16845;
      when 45 =>
        table_value := 17189;
      when 46 =>
        table_value := 17530;
      when 47 =>
        table_value := 17868;
      when 48 =>
        table_value := 18204;
      when 49 =>
        table_value := 18537;
      when 50 =>
        table_value := 18867;
      when 51 =>
        table_value := 19194;
      when 52 =>
        table_value := 19519;
      when 53 =>
        table_value := 19840;
      when 54 =>
        table_value := 20159;
      when 55 =>
        table_value := 20474;
      when 56 =>
        table_value := 20787;
      when 57 =>
        table_value := 21096;
      when 58 =>
        table_value := 21402;
      when 59 =>
        table_value := 21705;
      when 60 =>
        table_value := 22004;
      when 61 =>
        table_value := 22301;
      when 62 =>
        table_value := 22594;
      when 63 =>
        table_value := 22883;
      when 64 =>
        table_value := 23169;
      when 65 =>
        table_value := 23452;
      when 66 =>
        table_value := 23731;
      when 67 =>
        table_value := 24006;
      when 68 =>
        table_value := 24278;
      when 69 =>
        table_value := 24546;
      when 70 =>
        table_value := 24811;
      when 71 =>
        table_value := 25072;
      when 72 =>
        table_value := 25329;
      when 73 =>
        table_value := 25582;
      when 74 =>
        table_value := 25831;
      when 75 =>
        table_value := 26077;
      when 76 =>
        table_value := 26318;
      when 77 =>
        table_value := 26596;
      when 78 =>
        table_value := 26789;
      when 79 =>
        table_value := 27019;
      when 80 =>
        table_value := 27244;
      when 81 =>
        table_value := 27466;
      when 82 =>
        table_value := 27683;
      when 83 =>
        table_value := 27896;
      when 84 =>
        table_value := 28100;
      when 85 =>
        table_value := 28309;
      when 86 =>
        table_value := 28510;
      when 87 =>
        table_value := 28706;
      when 88 =>
        table_value := 28897;
      when 89 =>
        table_value := 29085;
      when 90 =>
        table_value := 29268;
      when 91 =>
        table_value := 29446;
      when 92 =>
        table_value := 29621;
      when 93 =>
        table_value := 29790;
      when 94 =>
        table_value := 29955;
      when 95 =>
        table_value := 30116;
      when 96 =>
        table_value := 30272;
      when 97 =>
        table_value := 30424;
      when 98 =>
        table_value := 30571;
      when 99 =>
        table_value := 30713;
      when 100 =>
        table_value := 30851;
      when 101 =>
        table_value := 30984;
      when 102 =>
        table_value := 31113;
      when 103 =>
        table_value := 31236;
      when 104 =>
        table_value := 31356;
      when 105 =>
        table_value := 31470;
      when 106 =>
        table_value := 31580;
      when 107 =>
        table_value := 31684;
      when 108 =>
        table_value := 31785;
      when 109 =>
        table_value := 31880;
      when 110 =>
        table_value := 31970;
      when 111 =>
        table_value := 32056;
      when 112 =>
        table_value := 32137;
      when 113 =>
        table_value := 32213;
      when 114 =>
        table_value := 32284;
      when 115 =>
        table_value := 32350;
      when 116 =>
        table_value := 32412;
      when 117 =>
        table_value := 32468;
      when 118 =>
        table_value := 32520;
      when 119 =>
        table_value := 32567;
      when 120 =>
        table_value := 32609;
      when 121 =>
        table_value := 32646;
      when 122 =>
        table_value := 32678;
      when 123 =>
        table_value := 32705;
      when 124 =>
        table_value := 32727;
      when 125 =>
        table_value := 32744;
      when 126 =>
        table_value := 32757;
      when 127 =>
        table_value := 32764;
    end case;
    return table_value;
  end;

end;

