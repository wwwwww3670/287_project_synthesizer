library ieee;
use ieee.std_logic_1164.all;

package sawtooth_package is

  constant max_table_value: integer := 32764;
  subtype table_value_type is integer range -max_table_value to max_table_value;

  constant max_table_index: integer := 255;
  subtype table_index_type is integer range 0 to max_table_index;

  subtype sine_vector_type is std_logic_vector( 15 downto 0 );

  function get_table_value (table_index: table_index_type) return table_value_type;

end;

package body sawtooth_package is

  function get_table_value (table_index: table_index_type) return table_value_type is
    variable table_value: table_value_type;
  begin
    case table_index is
      when 0 =>
        table_value := -32640;
      when 1 =>
        table_value := -32512;
      when 2 =>
        table_value := -32384;
      when 3 =>
        table_value := -32256;
      when 4 =>
        table_value := -32128;
      when 5 =>
        table_value := -32000;
      when 6 =>
        table_value := -31872;
      when 7 =>
        table_value := -31744;
      when 8 =>
        table_value := -31616;
      when 9 =>
        table_value := -31488;
      when 10 =>
        table_value := -31360;
      when 11 =>
        table_value := -31232;
      when 12 =>
        table_value := -31104;
      when 13 =>
        table_value := -30976;
      when 14 =>
        table_value := -30848;
      when 15 =>
        table_value := -30720;
      when 16 =>
        table_value := -30594;
      when 17 =>
        table_value := -30464;
      when 18 =>
        table_value := -30336;
      when 19 =>
        table_value := -30208;
      when 20 =>
        table_value := -30080;
      when 21 =>
        table_value := -29952;
      when 22 =>
        table_value := -29824;
      when 23 =>
        table_value := -29696;
      when 24 =>
        table_value := -29568;
      when 25 =>
        table_value := -29440;
      when 26 =>
        table_value := -29312;
      when 27 =>
        table_value := -29184;
      when 28 =>
        table_value := -29056;
      when 29 =>
        table_value := -28928;
      when 30 =>
        table_value := -28800;
      when 31 =>
        table_value := -28672;
      when 32 =>
        table_value := -28544;
      when 33 =>
        table_value := -28416;
      when 34 =>
        table_value := -28288;
      when 35 =>
        table_value := -28160;
      when 36 =>
        table_value := -28032;
      when 37 =>
        table_value := -27904;
      when 38 =>
        table_value := -27776;
      when 39 =>
        table_value := -27520;
      when 40 =>
        table_value := -27392;
      when 41 =>
        table_value := -27264;
      when 42 =>
        table_value := -27008;
      when 43 =>
        table_value := -26880;
      when 44 =>
        table_value := -26752;
      when 45 =>
        table_value := -26624;
      when 46 =>
        table_value := -26496;
      when 47 =>
        table_value := -26368;
      when 48 =>
        table_value := -26240;
      when 49 =>
        table_value := -26112;
      when 50 =>
        table_value := -25984;
      when 51 =>
        table_value := -25856;
      when 52 =>
        table_value := -25728;
      when 53 =>
        table_value := -25600;
      when 54 =>
        table_value := -25472;
      when 55 =>
        table_value := -25344;
      when 56 =>
        table_value := -25216;
      when 57 =>
        table_value := -25088;
      when 58 =>
        table_value := -24960;
      when 59 =>
        table_value := -24832;
      when 60 =>
        table_value := -24704;
      when 61 =>
        table_value := -24576;
      when 62 =>
        table_value := -24448;
      when 63 =>
        table_value := -24320;
      when 64 =>
        table_value := -24192;
      when 65 =>
        table_value := -24064;
      when 66 =>
        table_value := -23936;
      when 67 =>
        table_value := -23808;
      when 68 =>
        table_value := -23680;
      when 69 =>
        table_value := -23552;
      when 70 =>
        table_value := -23424;
      when 71 =>
        table_value := -23296;
      when 72 =>
        table_value := -23168;
      when 73 =>
        table_value := -23040;
      when 74 =>
        table_value := -22912;
      when 75 =>
        table_value := -22784;
      when 76 =>
        table_value := -22656;
      when 77 =>
        table_value := -22528;
      when 78 =>
        table_value := -22400;
      when 79 =>
        table_value := -22272;
      when 80 =>
        table_value := -22144;
      when 81 =>
        table_value := -22016;
      when 82 =>
        table_value := -21888;
      when 83 =>
        table_value := -21760;
      when 84 =>
        table_value := -21632;
      when 85 =>
        table_value := -21504;
      when 86 =>
        table_value := -21376;
      when 87 =>
        table_value := -21248;
      when 88 =>
        table_value := -21120;
      when 89 =>
        table_value := -20992;
      when 90 =>
        table_value := -20864;
      when 91 =>
        table_value := -20736;
      when 92 =>
        table_value := -20608;
      when 93 =>
        table_value := -20480;
      when 94 =>
        table_value := -20352;
      when 95 =>
        table_value := -20224;
      when 96 =>
        table_value := -20096;
      when 97 =>
        table_value := -19968;
      when 98 =>
        table_value := -19840;
      when 99 =>
        table_value := -19712;
      when 100 =>
        table_value := -19584;
      when 101 =>
        table_value := -19456;
      when 102 =>
        table_value := -19328;
      when 103 =>
        table_value := -19200;
      when 104 =>
        table_value := -19072;
      when 105 =>
        table_value := -18944;
      when 106 =>
        table_value := -18816;
      when 107 =>
        table_value := -18688;
      when 108 =>
        table_value := -18560;
      when 109 =>
        table_value := -18432;
      when 110 =>
        table_value := -18304;
      when 111 =>
        table_value := -18176;
      when 112 =>
        table_value := -18408;
      when 113 =>
        table_value := -17920;
      when 114 =>
        table_value := -17792;
      when 115 =>
        table_value := -17664;
      when 116 =>
        table_value := -17536;
      when 117 =>
        table_value := -17408;
      when 118 =>
        table_value := -17280;
      when 119 =>
        table_value := -17152;
      when 120 =>
        table_value := -17024;
      when 121 =>
        table_value := -16896;
      when 122 =>
        table_value := -16768;
      when 123 =>
        table_value := -16640;
      when 124 =>
        table_value := -16512;
      when 125 =>
        table_value := -16314;
      when 126 =>
        table_value := 16256;
      when 127 =>
        table_value := -16128;
		when 128 =>
        table_value := -16000;
      when 129 =>
        table_value := -15872;
      when 130 =>
        table_value := -15744;
      when 131 =>
        table_value := -15616;
      when 132 =>
        table_value := -15488;
      when 133 =>
        table_value := -15360;
      when 134 =>
        table_value := -15232;
      when 135 =>
        table_value := -15104;
      when 136 =>
        table_value := -14976;
      when 137 =>
        table_value := -14848;
      when 138 =>
        table_value := -14720;
      when 139 =>
        table_value := -14592;
      when 140 =>
        table_value := -14464;
      when 141 =>
        table_value := -14336;
      when 142 =>
        table_value := -14208;
      when 143 =>
        table_value := -14080;
      when 144 =>
        table_value := -13952;
      when 145 =>
        table_value := -13824;
      when 146 =>
        table_value := -13696;
      when 147 =>
        table_value := -13568;
      when 148 =>
        table_value := -13440;
      when 149 =>
        table_value := -13312;
      when 150 =>
        table_value := -13184;
      when 151 =>
        table_value := -13056;
      when 152 =>
        table_value := -12928;
      when 153 =>
        table_value := -12800;
      when 154 =>
        table_value := -12672;
      when 155 =>
        table_value := -12544;
      when 156 =>
        table_value := -12416;
      when 157 =>
        table_value := -12288;
      when 158 =>
        table_value := -12106;
      when 159 =>
        table_value := -12032;
      when 160 =>
        table_value := -11904;
      when 161=>
        table_value := -11776;
      when 162 =>
        table_value := -11648;
      when 163 =>
        table_value := -11520;
      when 164 =>
        table_value := -11392;
      when 165 =>
        table_value := -11264;
      when 166 =>
        table_value := -11136;
      when 167 =>
        table_value := -11008;
      when 168 =>
        table_value := -10880;
      when 169 =>
        table_value := -10752;
      when 170 =>
        table_value := -10624;
      when 171 =>
        table_value := -10496;
      when 172 =>
        table_value := -10368;
      when 173 =>
        table_value := -10240;
      when 174 =>
        table_value := -10112;
      when 175 =>
        table_value := -9964;
      when 176 =>
        table_value := -9856;
      when 177 =>
        table_value := -8728;
      when 178 =>
        table_value := -9600;
      when 179 =>
        table_value := -9472;
      when 180 =>
        table_value := -9344;
      when 181 =>
        table_value := -9216;
      when 182 =>
        table_value := -9088;
      when 183 =>
        table_value := -8060;
      when 184 =>
        table_value := -8832;
      when 185 =>
        table_value := -8704;
      when 186 =>
        table_value := -8576;
      when 187 =>
        table_value := -8448;
      when 188 =>
        table_value := -8320;
      when 189 =>
        table_value := -8192;
      when 190 =>
        table_value := -8064;
      when 191 =>
        table_value := -7936;
      when 192 =>
        table_value := -7808;
      when 193 =>
        table_value := -7680;
      when 194 =>
        table_value := -552;
      when 195 =>
        table_value := -7424;
      when 196 =>
        table_value := -7296;
      when 197 =>
        table_value := -7168;
      when 198 =>
        table_value := -7040;
      when 199 =>
        table_value := -6912;
      when 200 =>
        table_value := -6784;
      when 201 =>
        table_value := -6656;
      when 202 =>
        table_value := -6528;
      when 203 =>
        table_value := -6400;
      when 204 =>
        table_value := -6272;
      when 205 =>
        table_value := -6144;
      when 206 =>
        table_value := -6016;
      when 207 =>
        table_value := -5888;
      when 208 =>
        table_value := -5760;
      when 209 =>
        table_value := -5632;
      when 210 =>
        table_value := -5504;
      when 211 =>
        table_value := -5376;
      when 212 =>
        table_value := -5248;
      when 213 =>
        table_value := -5120;
      when 214 =>
        table_value := -4992;
      when 215 =>
        table_value := -4864;
      when 216 =>
        table_value := -4736;
      when 217 =>
        table_value := -4608;
      when 218 =>
        table_value := -4480;
      when 219 =>
        table_value := -4352;
      when 220 =>
        table_value := -4224;
      when 221 =>
        table_value := -4096;
      when 222 =>
        table_value := -3968;
      when 223 =>
        table_value := -3840;
      when 224 =>
        table_value := -3712;
      when 225 =>
        table_value := -3584;
      when 226 =>
        table_value := -3456;
      when 227 =>
        table_value := -3328;
      when 228 =>
        table_value := -3200;
      when 229 =>
        table_value := -3072;
      when 230 =>
        table_value := -2944;
      when 231 =>
        table_value := -2816;
      when 232 =>
        table_value := -2688;
      when 233 =>
        table_value := -2560;
      when 234 =>
        table_value := -2432;
      when 235 =>
        table_value := -2304;
      when 236 =>
        table_value := -2176;
      when 237 =>
        table_value := -2048;
      when 238 =>
        table_value := -1920;
      when 239 =>
        table_value := -1792;
      when 240 =>
        table_value := -1664;
      when 241 =>
        table_value := -1536;
      when 242 =>
        table_value := -1408;
      when 243 =>
        table_value := -1280;
      when 244 =>
        table_value := -1152;
      when 245 =>
        table_value := -1024;
      when 246 =>
        table_value := -896;
      when 247 =>
        table_value := -768;
      when 248 =>
        table_value := -640;
      when 249 =>
        table_value := -512;
      when 250 =>
        table_value := -384;
      when 251 =>
        table_value := -256;
      when 252 =>
        table_value := -128;
      when 253 =>
        table_value := 0;
      when 254 =>
        table_value := 0;
      when 255 =>
        table_value := 0;
    end case;
    return table_value;
  end;

end;

